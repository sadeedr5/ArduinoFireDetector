PK   �\XL�Q�  yj    cirkitFile.json�]ks�F��+,��n��/}��f��f�s�,�A�
EjAʏu�����(�@�gl�l�[��4z�@����ߪͪܶj�V��f��_�h1����]~��-�7�f�߮~k���G�{��p���UyUl��U�I!�X\Q ����AT�e�dz�R+�b��o�8��8������B2��0��^�l7j�_�Pa�T+�8�EɃ�(e�a��",je�p�M˄'�L�:�I �(�<��JD�1�4�+�\A���4�K�ɩl�9P�*&s�"�UB�@E`��́��V�A�d�}��Y ��#Bh�����$2�fA�)�!4z�&Ch�HM��,豚�YУ5B���k2�fA��d���C6B���l2�fH��S�c'B���N2�fA��d͂;��=v�!4z�$Ch��iA�lߩ6h�f=�)��f���f�AO�!�6�7"ǲ�Xv���ʎc�i���N`meǱ��*��.��ʎcٱ���NbmeǱ��*��.��ʎcٱU��]���ǲc�k�k;(;�e�V)�v)�vPvˎ�2��2���8��y�N�����3/ ��CW��\_pp�����3o?��WX~�ϼ��\i`�q0?��	l?p������̻2�����3o���WX~�ϼ��\y`�q0?�fl?p�������;a�fp��������l������3����C��@�� �\p������L��~��ˏ����������3�&`���,?�g:e���X~�������?��8���N�\`��g���<�Lz���.�3���o��1��gS��"\���,pYUU���|w��A��<�d��8Lڑ#�isN9zL9oA9�i;��S
qF!~��x�"�.R�*��P9w�i���O;�ϝړ|���n�s�������D���88w>�.A�?�?���D��z�ϝO�?����C�s�'v	%rvm�M
�!���a�I��M�����S^5�K�/xp_�ȏQ=�u��>�FM�Q#���Ӂ��M:�p��L���$	9�;��G)��mK�G�ú��O�'�� �����U�F ��x�0ꀲ2��H����J��U�F �� ��{Ѐa�@`���g���ڸ��!�:�Ø�	�QH��'R���	�9,|���gY N��a!��?sq�Eq�(��� (���q��(��&�,�XG!��ZA�`q\��8
�&����QH��k'X�8>�DW��v�
T[j�
�j��Q�v���Vc�X�'�
����R����pT�]}p�U\08�!���ꃫ�����io1hW\m��N{��@���j+�`,pڋG��W[5c��e8*Ю>�ڊ2��.�Q�v���V�e�~
.K����)���u��a���Tv���,1<,Ҷ~J//lB6xX�m��_^�:Dn�H��)���u��a���S�ya����"m����!���E��O9慭CT������[��i[?e��1<,�͂���[�Pi[?u��<,Ҷ�^����,<,Ҷ~�2/l�?xX�m��e^�:���H���˼�u��a���S�ya���"m�.���!6��E��O]慭C������l��E� (���KP�Y<_�h�MR�<�	(]O������@�o�<�"���������+V����	�=��}6A�3Т?A�3�?A�3�n>A��0^<�=�A Ƌ�>4�����x����L��m��;"L����Y/+���9���y:�+�@y6�+��t>2V�p��]Lc�m���cuj��j�j�<}Fc�g���������0�}�W I���ݷ����4I P_}@���J��WEF ��0������ �@@}	a�+R#P_�B���2&D�6.l��6�n�� �,vsX�F!U`8��7�p��!
�,�sXG!�`8�⸀�q����.��%�8.`q�tx������QH�'N�8.`q�tx&����Ǉ� �0h���0 �!	�F�quH Q�v���!	���S�F��W�$�V?)hW\�0X��hT�]}puH�@,`���Q�v���!	���C�F��W�$�V�(hW\�0X��hT�]}puH�@,`���Q�v���!	����\��
&��Srya뒄��"m���Sw�"+pX�m��^^غ$a�H��)���uI��a���S�ya뒄��"m����%	�E��O)慭K����r�[�$i[?%��.I8,Ҷ~�2/l]�0pX�?u��.I8,Ҷ~�2/l]�0pX�m=��S��"+pX�m��e^غ$a�H���˼�uI��a���S�ya뒄��"m�.���%	�E��O]慭K������[�$i[?u�(�$a�(��$a�(��$a�(=�$a�(}�$a�(��S$a 0��l�$ ��C_GM���`|x賡)�0������i�H� `0^<���I Ƌ����"	��xq����Y/-	CG�pyvA�����<��FK��Q�]L�%a�D-	CGy�_FK��Q����B���~Un��v�T��<\��5�ڭn�y��U�Ym�J��ׯ	ɡ��d,u^��E �*
�Lʠ�y$´P���%x��~���QG�CG5[���9��G�"�A9xD98?=�eJ�H<��(5!��Kld�8��ٔ��rd��IG�x���e#��_�����H�,��	-!��F&�_���K\߿��e3��޾��L��\��kMS���K���Yԓ>G2E� =��s��V�ztű�{9|�,�jN�C��5�<5�������Ya:��������06����H����g�@&@�D����`4�2�Ge2�a�,K��g)�����<al���9���C���BJ���ˇ������h��6@Y|E�t�}�
��o|!� C�3D�=�!VT�N����Y�!�> "2D�GDdA�����,�}���E�b�`����!�H^���.*2ơ5��T9 ��1�iT������qh��� W��t�C�5=�W�t�C� � �
@<�c��< �T �)��&I���O��FM*@<�xjc ��qx�W1$<�6�ϡ{�Ã��ϡrM<_�y�~X~5k��Z��� ���s�V��������C��x����8<����*���>X��A���P�&���Q:b?,?��4�|��qx�a�9ԣ��k}\�Ã��ϡM�w����L�x�%��K��!�A�!��2cCt)f��ubl�.G�]��@@��%	��K���!�,3t�116D�&`�.�e  Ɔ���Х���]���t�����0C�^2�]���t�����0C��1cC�+t�b+16D�)`�.=c  Ɔ�:�Х[��]���􉁀��0C�1cCt�f��bl��S�]��@@��u�3'�S�[��4�)��bi�l�	��Ȇ��؆�|Yo�FN�>�C���jM�"'L�:�����`�Շ<E0�`u�N	&X��S��IA��v��` ���)��$ �'���S$~O�F�x����r��i�����wB��e���p�s��b�㒋Ѫ��K��j�<n�������8�Ѫ�'lR����'p��?�4��y��;#�0f5�/^ύ�/���4e��F)�hefL7Ќ�f(7c���hn�s3��	��f���af3C���f�03����Q���q���1�7��'�qQ��eA�a KY�`2P�����J/���z{���e\!�ց����$+b��#���<�U�%��d�P<*��2/���G�U���.K&4f]���z��E�VU\F��2�q-k��R�
�T[�H'�,3e,�F��m�"�7���[�����PB-���܀lJ���q��}2���|f	b;��PU���K C*��(7�ϣ�k��	l�U�noD��y��&�ّn����+a/�n��w��.f��]��%���+:��]�aWln��z�:
%ͦޮ��no,=*���÷_�[�J�����J��і4\�U�7W�K�����+���h�M/��j���2�뛍��x���n�6�ߴ7�����]����[���:s���v�h�s������O�w~Q���;w����5�Z�okտn���C��<��7�u^�o[#Q<L�x��^��DS���}��vx�|)�͹�i�c�smYC���ӱ��$�$�X�H�W"�^R�ޒD���Y�į��uG⋹N1����F%����m4J޳����-��p�_��XF�0��,^�I����a�dۥ8�m�NN[������z�=KN��#⏑һ�"qo�㣁�{|�R}62[�E��="�Ή�ăs��9��ɇ�H18G����9̺r�Q�3ʾڮa��w��<�9���(�K��,��Gu�2�&�Ģޮ+�.>^v��r~q9�������|q9o�nK-uҒ�EP�\.i�i�ˉ�	e�����x��f��������YYd����s]��B u�c��q�<�B��5�?�'�лE^gz^Zy�������U�Eur?�����h�,�2����r��ݧ̂��Ur��z_��?�������Q���.�>�ɋ�f]#'��uR�L��]t�W�Q��f��QT&�cS���v���Fm�P
V�*�f��1�D�'Ou���,+��<r��Xow�M��;��q+���uy]"e)E�������7��Rf��?�m!�������*6�a�E�����l����q�%�{^n��ߪ�U��aߧ�^_"Z��Z9�k���,��H(�Vq���DyN��8J�y^9XR�R�J�/
�eRyf��\���)/k�r��L�����?��rV�Yt�<�Pa����B�����vQ)=��XzN�TYU����������mS�vj{��>^^nf�o�����>lo�~�̌�]�V-f���̶�{�G������ۭ�:o6�Vݨ|����c���+�V�s����[����?&k~�T~�ǁG��n�7�W�۪��gs���a�#�{��p�.��E��K��$��cy��d��y��B�:�H�j�(s�e\T��/rg�"N�QO�N�.Q=�`8�R3�9�|�(�æ�-#}����-I�:�N��-=�d�L[;�A=� �#���pt@{ �
��-5��+1��e��Ǘ�T�aV�E�Km�M�TqP�K.�PdѨ4t�s�Q��O8��3>I��=Qzr�}ؓ�,�IƝ��Z~�θ�Pb�l���0��Z���R�ݶ}ToX%�]{��a�7��h��H���U��-����yqw)_6�?�����cBм���k��������z s:��쿩���O�a�O7y���]�u�$�y�0��a���Å'a��f����r���|��<�6�tD텾�4���C�{��I����Y�o��H"��G"6[x����Q4�Q*bY�$I�@�nH}sb^繮�b��Qa`�S���϶V�e���i	���}Ҿ�Uj�⟫��$�����^���U,B����V�T�,��JG�1��V���^�tv�V�_�|��n����~~?�v����_���-c��.�/�l�L.uv��4,N�<�u�H1��zY���^E���}��'����+��j�g����_i�pK��8�t)�,�2�e��q�e�����V����3���V���W�:9��Rg�I��	p�Љp��R��ٰd���9�W��>�[{�ݺ�o��σX,�"h�l^��45��j��eI�)MÕj~�2�(����d�Gئ1/�T��}���V��~mԻ��ޯ��h��k����a��B��Z��6�G�.��]¦r����A���Wϲv�E���ש�w����l���U�����rnz6~�_�����3[/^�?cy�ru�wp͏�p���9�{?�0�NF��t9����q�q�>%�(gP%:Jrz�zGI&�
#����8g��\���C	�%�%�9�n7�5�)�����Gq(�ӡ8ԡ8��b�=�����W�g�P��0;��(��Q����h�K%���dT���pʨ��їt�q�xul~$���|2=���uߪ�����A�6p��+�'}���<p!%}�O&QC�t�gt!�)����5*s�2��g�D�<�B:��9Fv����h�1�ۚ���G���I��8G^r೗g����.�����%w�)&�{��w�#/����p�\d���P��@�̋nݨ�id�L�d�98w�U�|.�I��sF�p7��L��\須�I���SZ�m�٣\ȼ�h����j�|mTѴW�_����|s����^��W����o>�?�PK   �\XH�8�  �  /   images/273c8146-c058-4dd4-bed5-b60da603675f.png��PNG

   IHDR   �  {   ���  JPLTE   ���AAA\Z7��� b҆�� @P��V�zӃ��q�������♕b=��V�R{� .Z I~z� &h��f����..1������"��G�hhh?{� `��������� 2iUUV ~�nu�  ���&&&��󡡡Di�`���m���)H[�n�q�����b`^S����e�;6/BnmmFB����� (C���:bj��_�  ztm v�3{�/1%*_�9998L�5Z��㙝� >ry����f5Olvtu]u�~�����  Jw�$?|no���{|N|�ς}vp���� ���y�� 4r    (H��DN�   	pHYs  �  ��+  ZIDATx���_����s.��p(JdA.j�]&��u��
�S%�-�!�����E�o�K�VO�I$=�����{��I>	�C���;S쎏���'�xscR`2ֿ���C! ���)��iK�;&���-d(�y!I&����BF�1ż�&c�P�n�R�t~�Ea��@1?B�(�bl ���l
A��N��@���xSl
d>g�,"��)�(s�X�D!�qN��l�}��"��x�Q�f��w����(�3R�z�|(x�|(�K
Wxþ|(x]8E��L�>��A1YR��YR<0
ޘ��()J����()J�?.E������()J����}Y�޳�_*E��Z�"�3�|g�R�;�� (&�f��<�	���ϋ��c�%��bҕ��+++�����$��=�&�+ow��s��1
����z�Y/)J��C��#w�P�6���)~�v�C���s�M��B�W�x�C?��s�4?��-�8{�Q �SJ��*�|)��R��ٙ���1�
WggW=�X�5a��:0�������j�{�}^��1��ulW�uF)�S�Nf^h�(�U�]�y�2�B�^Q�4�Z.,����^�.��XM�غv���0����t���S6�Q�^G����0J���?)B�G�f��o�v��P���q(j��ԭ=��]���ا�����'J���H�\
>
�@�{o�Vf����5)E�;f�^�Q��:��T^û�oR�Pw�>2�4� ,���}��پC�O�Bb=�2�N(^w�(����9���/,�����>\�MA�+t����~^d�1�XMj���B�Y_N��&�=��
����VՓZmJ���(���A��/̸֍G�Ngff�R#���v�N�x���'�K[���Hjg�Ç���q���z������/���=�)�W�������o�ݒ�{������}$*w�r��?�������h$��e�3EF))J��(��-FIA�49%9{^�kGEjƉa'x`̘Dkx�mg�R)�a�Hv
�bC�Dyk$Q4�J ��W� N�1 �9"C��a�>�g�L �&Ku��p:�P
����F�����zIVc���xC�Y*��.P[����4,	@ qV��N
K�6*jh�!�B$�a�8e*��KPx�l[TmK�s$*�����h�6@�� ���(�)�Ԉv� $�UL��c�\��h �)x���uS�$lm��&z!Q� �'8�!�tD��=�xD���D
zt��N�,$�g�E�LUEl[�X�0D�Q�2I��
B8�s�E	l��"�� ���Mn��*����MS��-pG�h�-��m۾$|�&�B�%�}&���񵟈�S�bM�@Ѡ���|�J�BP�/7 D_ =*���XM<���O(�a��H�B��ܫ�1&$�7�PX&��3q7��J�	i�ݨ3�BAڤM�\
�����;�����*m��0pm!A֌�I��	i�(��t)NDwOJQs)D��$�.w٥#S�&�r��4��)�G�5|^��?&���4�m{�ְ1e˒Q����u�j�(�U�PA۲N��a�fYFQgfX�L�*;w��)��eH��K� �2�������:i���s�Ƚx��l�� �q��VI��]���N���U}��S�(V��Q��n�T�ˇ�哠aR(`��9̤IQ]&'J��7���M�*}Gz�QTB~��d�amq?#�E�����4ۅ_s�.�=2���	Q<u�p%�|�RXveLhe�E���
&��'UK��'����S��WG~	Q|����).K����()B�$D����ɿy(�:�4D�iC{~@Y����")��Bϧ	�"�L�df��%�`�"����S ����s�'���"TT2E������-�(*R��ݯK���GƂ/�6�"�a��~���M�����cW��5Os~wo��	9��~�kDM���X��K��fT�~o�Q���Ƨ��̢�%��Q��͸>8b
�H�M���'�=�2����Ύ��wiA�v^��f��������ut�%��VG`�x
{օ�|��t�N)�}{UW?���u�u^
�F�K����Q�#OFm��/n��G�X#Po��ka���n_���"���Z�����N�r���-�ԑSl�S���B/)����+����R9,ES��ɿ��[��~t:Q,Ew���b�.|bg�[,�}ݷG�����]z��\(�ۅ�gK��~}���	��D�݉Sj���[�}��Aؼk��������/u#����ۛ�^ݣ�x�j'�?���|es��@,o^�zR$�i1��ʦ����2yx�l����B(p��.�Օ@�޴!0�����­�q�i�����������A!&�0�+�kM�.Z�1)�!1ʋB[��l����S�:�����]E�bx����8� rv�p�(��NqKo�q<�2]
b��T]T�plQ�mq�؂ګ(��A���.�e�}}�a�J1�̃��qZ߯F1qt��7i����+��~ߒ�������Ǒ��G�;�#G�r�^|"c�a`츖��
���5��|os�s�6W���O����#�4�^���h��6|R�8Ɯ~�j�x����ณ8��3��m+>�]��c9�~<����[�q�X
P�B�%��}oVp����O-�bbg¥p�ً���6��wV�ΘV �����������nQ�H�.�̽g���������Q�L�j�w��F�U,y��R�ӷ$�B�|�p�~�b��K�ݼ�@��[|d�<�P��)��L�������#�,���ȓ/�\�}?�a~�)�tQ�D�)�t�t9��G�(���f\�t).r|������G)�rpp}}p �g��d�� �g���D���U��2���V��2#�P��b��U�^5�흃⥤�N�F~B���5*��i�) ��8�7@Jb>[����D��o´��{�C����E�!�K=t��@
��
�_oT�,}��X�� (�->[|.m�l�,k$[d�Za�g�G���]�IF����)�w��ol��Џ���ެ�{����s,o����G3H�{�杓��=_#r�EոaY͸�j|Z�9lq'�1Qi�Q�%��!g��{� �j(�ij�!�v�7G�Hu���+��x%i> Ek˕˭8���g��V˝
i�W�0����[1��j�9:��ι��s1 Bec�Ξ�Qs�1_|a�Zl�-B�b�ĭ����r�PP��Z����)��)�!&H-���bq��H2�(��~�x�q�i��W�3��&&Jd�K�#ڋ�lO���r����S(�J8+l�J��jy��|_��5��
!��s������l�9@TB1E"9u|M��i	΂I�e�����RE$��l��Q�Fn�H�#Z���d4�LapRo=vXg"q��څ�6*����Gq�i������D=���nE����9m1��<�%�������Q��ϼ����ѧ��"����F|���r��l�f9-�����bN#�c��/Q��5��� ��-6��Z�fe�x<Z[����c�L�7��޸��X�S���@A�aY'm��E���Sol��k��!��K�&R���]&<��@ݗ<��Sm1Z����a������GQ�£�lA{6�I�$�$���y>�V�F�O9_,Bz`��, N��4����.� $j�|;&L�U2���35M#+����25s
�Ml"��C��)��!K�O��1����i�V)���VC��P58��HfY����(mQA�� ����\3h����+�3�b��R*4�@ 3p���8OL��L�SI$��U�5ɘb
A����T&�����B�#����lJH� .�_�*]�^$l�t4�z���)pE��::a�:H��F��>��� �P͠W�~?�����)pU9˔Ԝ �P���)��۵��kEk���� �<*���LԶ 0��Qcz`��42I�聲R(�eྦ��l�P�RM�.��]�*�%� d��1�V�Y
"�|VA&%�"���Ռ�(�بm�����MD�f�7!w`ȸA�+h�7]�A:���Z��p��(ȗ#t��P$�u�QH�3��!<<n
`� #E�$:u�I��1�2�%S�_HR�YҤ%J��9Ȏ�n6��������{w0�NP��a"�zx�D�Լ�Q5�����U ��(��Z&��*���c��P,bY��p5�e����I�� ��X
W��� ���!�C���HQ�bc��m���P|�=��n�5Rd���-���h��Rg�������I�������~���j�3x�7H����JqL��E�:K��E4ߑ��#���d�����h^��FW_Ulh$�O��.�RĽi�S���R�)�O�G_w�A=~��2(@HXY7��DE��R�Y��0���O������dKr��_I���P�X��ic>�8�7���$M�*VsEʊ�����DI�h�%EIQR�%EIQR�%EIQR�Y�(�KQ%P`�b�.�f��x�K�(VJ
OJ
OJ
O��(dD���    IEND�B`�PK   �\X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   �\X|�K�?  :  /   images/54ba0d46-ef45-4902-8525-adba90967d59.png:��PNG

   IHDR   d   9   ��}   	pHYs  �
  �
܄߉   tEXtSoftware www.inkscape.org��<  �IDATx��\il\�u�ޛ�f�pI����Z�Ց-ٖ�ڲc���I�K\$�Q4��-P (P)P�E�.H
4HlÒ�8v$E�,ʶlY%R�(R�D�����3o�9��g�!9o$[4���{��w�=�|�|��G{~d�KY2�`��)�� �"����P��uݪKƒ�%���̝D`j
��~�u7�I�M�]*�2:;��D�����ї�R��B� *J�v������4N�oCGo�f����.	�ޭ�Kg14>�OT�3^���
)XZ�1�z�U<�3�U�iE����3qT#�V�tb"���,i�D�&.�������E*b�|0��I��	`p���,a]�pg��!����BtC`�m�6`7V����-C�if*�c�bb�\���z!MHhp"�r��H�{��
����� �*��5tNQ0c`�5�^�ċ�P�1(�˚���<-�t��@M׈�;VF�,e,Eq�
^��?��%�y��D�k�aM��i$����JSt�a�2|�q��Pmx���g"״ӿ�[N}��Σ�|k�RL�cMn����4a�]#
&�2�ۥ�R���Il�I�aEg���5�����2^��C���t�{"2�aG.��ae�A��!fϞ��XQ�c�k?�3�}.���g�
�4X&�NI�K�"J���b��t��&�R��;��G�K��v%-�[L��P\�ώ�νF�RV�㟞���������t����`��l&���S��b��!c��)'��<�9H�:����;;�
��'��	���4u"m���������h)OQ-�M��5���^X��*h����Z�[�YL��W9��j�*�P�q�
9jŋ��s�b��l�bN*�P���7N�|�iK'�,^�1�YH�ѻF3c�]1|go[v~k��Bow+j�ޥA�q�ݛ2+I��Ԁ�m�aˎ��E��wI$��#<��KU8N�#]�9�I�jX���vʹ��>�{<fj�2L�<�T�M��dv�h�&H��#A�UB
��۾��i���m�e!`\��cmu�۰������u��`o�E���dn2)ꩨ���_�.� ��mD<Dc�{��U�����=8v��(�g���}^Ϻ�$+������+gttk��ɻ�\��
	M"�c�c��ဒ�����9U&XpzsnR]^���,M{?v|N�PFZ\��T����/?�!1N��D�gRn�E��aB��5'0��"�N�yv34��{���d+ *�
*�3��i�΢���ue؋{z�q����6����7��y����Q���KN`3����ښOBv(�TB�+|��~7�d\�"�o!(2#�))��)!���V�M:B�UJ�	K�-
�П㤐�A5g`�tT��,q@�u첏½ E]����Hn�8r�,ǩ�Se3=�._8�D<J���KU��S�h�&0:m@^D��������*=+
ajj
	� �{4�SGhU�&�I�y�J1S�W'�8lB�h��ب����k���d�v$PS��ehtZ���M������TX���xh@�H�D
�)�G���ĉ>����-��b�ڵ��|���J�m###���C  N!���*z&4L�;���x�xf}?�]+GW�WX�<O��t�_<�]��?���-C(6���BD�d+z����eӕ?�BǗz\�4__�p_�B��HsS��-���|�rlڴ	cccp��ęFQWW'��-f:0E>����m"�Ǉ8�k�o`���	VJ���4�cI+�݄D�mu,�E�ɑ?�(�cm+��Qz0�6\;�{���t�Đ����-�ᩦ�===())���J�Omm-��$�_��r"�_���˧u#Fn�Iq����G��c]d!㷰B��B>�S�ô���+u���"��-�
��;~f��RyL3S�笨��*�"VIȄ˲}Lf��>�-��y,���-��iݺu`ٲe���Fii)z{{��S��W>�ah�1�-4G����:L��2�[˳1�0?�KY!�,�{�yrg�oI3u�1�ߵ��H�ȯ���g
gz�Ǉ��Jh��h���,� EF��Cn��C��P[+#�e�	����x�^7^=��gs���0}��[��h2n�K�� '+�n�O�v�s_F!Iz���d_�w<�zb�}�m�L]�i�N�6�H�{Las�^��� Ɖ��6����k�<(X�a�G[��[��G���J�N�P������V�s��w%�򦞇4��xd�"���a1��N}�2<ͮ0q�0�g�:���uS��o��u+7 4=�}��?H3u*�wm��=�"89�r1�X_:�7^�g��w�OQ֓;��`�|�H~�4MDSl�7o�������8�����ֆ������7���12�+�N�^�"9|�Sز�A���Ng.?���(�k��.�6��dX�]��,n� SO9z�B�Zue��ML��
�Z*k�aG����QgX!l!�HD(�C_�׋���crr��� _f��=A�\��S�jJ�������8�C!Y
�����"|(#���f��1����꼈�k�S�L�cS�<��##=hnj�0��m'qc܃��l��pꜹ�G=@/����[�X0!/��8����Nu�YHj���6b��~�r��5�1�:������
���_i{l'��'����c����'���^���:5��76TkH$����ԯ�8t��^��!S�C^?�6�/�J�I��V�&Z���QL�y��8m�AUd'u݄�2�IHM�9c�sb9�\1���}1���
�Y+���0��j�I���py`Sg���i	)�E&ON4�x(*���[&�$|�a7���/~)���+�[<��':El���Ԭ�v;��/��,`�R��U2q�����~~<���P�c*Z����J-h�YU���c��D	q�x<�Br�z�L�%��ڐ��3�d��������D�NP�rT"��f��g�)+�7�o�:E<$�ȋ�iO�_���}x�)k開9R���W��/�"�W�`[(J��
��y	eqL}v9��CK	��pTGRـ{w,�A┄�R�L�a�(��b�R9��K�	�:�6��J��On(�����GX�@#���rV�
�#N�i{��	P1L1�ojM=�ZS�����L=.c2$�f�	�&Tl��A���B1I�[�DV8I�W]*�NqD�˶�C:]j���F!�n-"i��<^�9_�P��!���{�o��E�4�#�p�e�S��1�ƎSϾ�"��cxv���cYL]��Գ�f���L��HX���������:I8�lI�5�ۚ�輢[V$���"��41,P1l����f���~/3����w>������ԯ�2���'��u/6m���k�ޡN�d�y���b�|F8�L�*��ܚ�+�HQ�dV��n��C�h/�:�HHs�a����k�k2L}3��(9 b�W�0��-�^��.b�!�L�s�8�S�۶4�c�T�d�آVYsNx��2w�|9�n_�L�o��ϑ��\ԁ�ky���p4[T�$�ߖ���`u����~op	Υ���L����i����2�vb���[.���b����=���S��@r@�_CE�,L���
c��7e�}C�K98����:��U�~�>`ny�,}o�v���כ|8�❻�A�v��L}������Ś�ś
��2�O���$I�Sk�t�8h���Z&�ԉ))�F��b%�����u�H-E��l`r�?���@�8��+�x�`΂X���y)�����G�ig.o����b�gM�Zs}�\��X���kK����<�� ���_>�)�����^b�.��6�:��{\ؾ��
Νw���Ҏ0Qt����M~�+6̵�����9#��w�s
���8#���:�S��[T�� /\�A�"��n,%.d�s8�o���^��=��lhY����cSm��0��8��s��FL�� ��E,�k�H�N��hO�����
�Iۻ6D5)��k����pb([eN�����VT#��V	�,�ld���2����sp��㗼�-���n���`.>����d�G��3	9�MvE�[{��1�$�^-��١~����nii��ѩ�HVf���Q����1�ӓB^�3\\)��"8��L�ڶ�Bǲ���&��
�YS������r03���T�����yI�^���C8���ؾm+zk�7�n=�!3�%�
L|g_m��V��"_署�?B��<@L=7��N
#-<'��`�x�dQ���{��j�$|�7���~�%���f�S@�8�ѹ���9�Z[�DK�V�VcR�?�y����~dsO�J`��oaͺ����7��Fp�_IH�);&���cϓغ}?����q�PTVp��`�W�m��ԛ��X�N�!��$��N�ʀ�s׵y�է	��Gb�w����̄�7{?+�0uw�
ce���y���bY�����38�:��L�骚����s�wiy5��F�޻o� �4N� �b�ǋZa�g���c�<r{�����L��X�ײ=���X�ǩ��Ia�l�h:wDN�M��H���oR�
�n��Ŕ+:�t���5��~�!��r�k��@_O�`�-�^�ev����SoaA��X?Z/6����b�|/f���L�$9L����
���� K��u������|A�;/�?�+-�?I�ra�����v���:AVbDFd
E�o�{��8 {���.�z��R|xqQ�9�X������N�q�Y�������ݬ���s*�e�M]�+]N�r�h0c�Wۨ�{�؞r�盜x��4d�W<A�����Z���ɩ�{��EE������4�Cq1��7�xL�9���|�}�W�'/����mI4u[L}z Y�Sg���GW	3u�a_T�Rbq��è_^v[^�dK9r�*Z�F�BBv��SwQ(������a�_>�tSN�1�����0@��TZ��a�t1E�xvb9u�L'jȖ��}t��Р����z�O���d�c��~��_xɉ+n+�o=�sj�۝ضJk �T��^�S�T��Z7�e1���%���2�n�⭋>띚Y��;�j�o�x�rRXH|$U�)l�7�"J� �Й_T0u�2���\Ԯ��"���;(�_�	5���(w�,j	�{�6���k�/�.Y�mw��e�#�Ǩg�-T�^��b���r_��UYb
�R�8�WKڞ    IEND�B`�PK   �\X��@��  ֈ  /   images/6b718467-4333-41a0-af30-09c4429f5121.png̺W\SO�5TD� �H��A� �7�E:��((Ho�BCoI�U��N�H3��	Ύ��]��s�[6��33�Y�Z3��kM%*rFrD���R��	]yq�:pGWwwx��l����,~D}n2x+y뺿���������9�9{�X{��{�g�I3�@�A*/���g�,xd��NG'���z�Q�H>��?�`NT��(H���`(�w>v���Eꝭ!���h���3O��(N��k�Wcclq/2� ,)Q�̪��t��'���M���k���x�_�Ҍ��9�#ūW �G͔���b񟼁D���w���W�/V׼���FM|��o������俿��˓_;����wcD�����i����F�x����mR�-C�T[�,G���Fn�7Ū����=1Wð��pm�~����Yj*�-���ҩw�X������{F8h.ӹ�}o���)�q>m�YG��G���5�J���W~�uP�|�_�_~Pf�)���?=M����"P�ی���C&�ѩ�ӽ�M}M׀f+~�ߞF�y>(�<^&V��==����fΈ\��Rd=8�h�2������W�/H��X��g�{;!��h��=��X�H\��QZC�Pӿ��o��i�:]�3	X�|��x��q�	h����#�.��nl��ںY��ۤ�Og)hF$��� �/TJ�v��Gf�����rq�vJ�R�y�I`���3�*�z=5�+Yͯ7�I��L�sD1z�Ё�������� ��k��Co�����M�����ޫņ���8Ϭ�����ps$�_w<&j��4[�J���f�j^�5��]\�`�:jȚ��j�7�}�t��2���JC�ܖuڏ�vEOO����O\�`le#D�5��s:iͩ*֮9+�q�37�d6A�U��cMG50��Ȣ��r+�9r�~?횓i��U�H�G'ŦW:J�~�ˌ3�2� Ο��}j���	~Y���?\͘��V,B-,��u��FI�k;��ޞ?/���hz��F̃�ŉ��!��w%5(�FI��� ����`8�  �j霡)/�Nsi3O
}�!��k�̉d�b�
a1��t7����*"(@��	3����	��6e��}�X���t)��V1cq�e;��I�	�A�<#����\����Ĵ�V5y/r�)�l�/7��+D����cPf�e�g��f�YO��]�5 ��ΠjO��U��7�y[ň�
h\�T&s�]���-��Z,�WR��$w�HA�O)����"���Јԍ�+��"��`��z����U�9;#f3�Ĉ#�&X7��|�%H)�77�#����<NA��\�7���O/��6Ź�L�2�CFBT���;�G�;����4�O����������;[B��N��ݵP.�wJ�r0�z�ݸq������|����3w��@���a�-(>�]������������2/��h�����_���]B��Z/2g����@����ۤ�-����A�	<n��}b
�2���i�؟3)��]3�>�>:�b��Ky���($~�-,�dv�%�ğf���l����GT���@�����;L��@���b��x�mp�[<5Ե�US���H�3�ִҮ#�ڗ�,3����w+�kT,Ѷ�x�Ia�h�=�l���7�Q-nTZr��_ߝ���)�i+Q+���E�v}$�g��\6��1����[d@���c�'�w�3���4��3�K��<Q��C�iD��&kel�;Wh&X���8x��Yi��k*K�����껅�5��\��!���ٔM���y"f�&俩���Q�5b�e3��b����X��/�~?l�	�~Q����{�+���5��'%��E�)�|����Fb$K��>"���}��~�3j��i8����속i?��"�k?���Z#dވ�)�]�`odևX�خO�����L�r��d��1���?��m��q� ��0]����W3�[�����7M��Q�����\�\�w;'4%Wƙ�h�O`=e���Z6/C��ݨ��H����g!���W��� ?���}|���ܼ��BpS�z�4ҸEmF�ٯ{V����7���I�4k,4T*����B;��z�B��Ɩ��D|9j�:�q�������������ҳ�D�&�/6��^��I��m�B�,K�͋igd`x{6-'sj?��u���5�*]�o�YH��,���6Z��Lz<�Ŧ�x���WJ2<nB�,i<���^+�WJK<n<�L)<mǳ2��An�,���q!��o�Б�u�Wk�Ğ�r
����>�01���w�x�?}�E^��A�+�V�m�臹b��LRP�I��<��+�'sؗ�љ/z�0N}�&�4�P�e�(��x΅���Er�Y&Hڡ�6w#��n���a�����zv�K'��˕v����̩�����sE'ה�?>
�9��&�!�O��vL�-#�M�R��+�������zm�\qBH���)o��v]jv-Q�!+V{TΖ�J�z9A.�����E���Edܨ�-\��*��q�M�O�W�F�0���C�Q]̚-���B$��������L`�!.}Y�4M>5�
Zb�Ub������V�>�s.�)Lx	W@��h����Vϰ�&P��z�������Rʷ���U��q�Z��kf��k���F��{�T55W��OL��9m�������H5�η�-]J�.�t�D�@���ݪ�9q�c1G��X�n��t�BO�79 �a0DW�e��+V�#���s|���c[5q/�@n=�ŇؽP���p�P���E�b$�%�1Č�lo�QHN/h'��8t���D<��a�]�dP)H���넆�}���������h��, ��0jaη؜�����ԡ#�҇-R��c����ojFBs�9����R�ֶ��NڤubA�rw~�Py��l�N�	��v�a�{>9���X\՗A�[�@�����}#U\_�+�4�,����7[�"#�Rv
Ȧ����⋭q�.��p�ϑ�Jz��c�Ve?������R&ΰ���I��\��cc�?]�ș+CW�`系W�����������Kf�_i��S�I�K!*\��"y��U�篂(:I��d~�V|��?�>s���'�V�g��<��w�ش��CH����߂I���`���-�Xe���,�'U�F��8�鶵��*`1�d�z�����rg,ǁ��\���d6N��A���Y��<��WA;��-��4�������C��rLӌ~k,0]���{��U BÚ����z��m]#䐐�I1K�$�����k��m�
}�sgɳ��ug�Sn�R�/e�?EQ_=W�.�+NC��_�)���q�lf�F]���Ms���(d�2|B�q�A[��6��(X�����'~RL�Z%��D�h|pg�� Ձ�>�z�x�+��n^BB��0Zᐂ�)�����؜CΫ���X�rK�dA_�R�aa�c~nT#c��dD��P��w5��m�!�T�!;��	iN��
W���陘���4M�W�N�sq�{���f	̊�d� U����Y�_�������~ST3V�]�?�ŔE	i`d�]���և���'ǜ�:�f���;�nqԬ�f�O�r�V��L��A8>*:�0fV9�v�B��8�P�w��wXc�4��N�ڵ��>���ֳ�n��_�������ɨ���i���� ��.:��꒖g�$����(h��~&隕���w�am���^�j�9I(�8�>N��L[�6W����΅2|(����ܦ��Wo��K��LH
6��q�I\�x�X�DM҉�<�'�mk�wmC��-U{�|�.�:���z�E��L����~߿μ+��u�����]�7��xQ���DF�r	�4ҞV�j��!.�P�8������Ӡ/�?���w�PҮ ��ݳ\zC�}C�ܵnË�iMY'�8F5=��OU��� ~�v�FN�3pl�<�����,6%��!�X?���+�D��P�VC֚[�w!�<�L���hTg*v�X�k>��m�2�:ɏ��a��K���ƮT�{C��h�:1QY�=3m�i�o��e�m���'�v�Bb>� )Ҧ��`%�z�N��3���hXO챟1�f���R\��Ԇ���,�g��3��W���j)Z�В��ԑ2hʆEYc�et��VE�j�!k���oIsO�lU��W�j��~��^�t�D}����@GĬ�����������,�}j>�4�w
��>jvNyY8ug20��ڳ*'�=�VC�ưۍL*�Z�F@�<~��3���N)�pRص��G��m1�
�a�M'ud����[{�M���"c�V6MB�ɓ�l�P�L?����?�Gϰ�<!����e$K�	\D"c�h�8?�q~:H�qq��0��I��Tʊ���|�@�+ 獸����@�`u]���:o��"��ݚI��;l����V��	5R0�}�i�}�(M�4��wΖgN��l�An��Jq�6�7�V�^N���j�&�����\�A|p�~i-~RV�Z�m��uMriiQ�u�Xd�d�����ː�$��A�$�����ee��V�W̌;�A{Y1�D�8~y�{�N����c��1����M02S��6LquW�6vbΪ�5e��`7[ �إ��?�*�t�$�j�D������'�Ӆ%Gxc5tz���kN������Ͷ:�xxX�9�Ji�O����c�d��g�UM�ٰ{�ro!,0��n��iB/y$Bj��v�hx�v�wz�(��?ג\^������qf��u��j��l�׎ ���"A�l`��aߐ�󥯠��w7`��%-�V0/�����o롦%-��΄$���#�B ��Ŷ����r������q�S�T;yJ��ͯ������>,��*M�op�T�צ%��CM�&׌+Hw��n2�.��9��~��$�I�Z�ʋi(��Ғ-.[�mj���6n���T��Kb�V���m!���}T��CM%؇�9�||[�������Im�2C��r�H'?�9Ƨ�'՚z���۸%a�rK,�4�_`&���d��~ߏ8^�
�_�"D��������3L|+Na�SL�K
ł��b�U��|�l��A�'G�Jq/j"�0�L��i�	��B-Jo0�Z)�x��έ��S���������Vם�,���ON�>����h��X�.��4&�Lg�a�f	T�0������I��Y�E�t�v��8��v$!����-�ᅲФ���0zyj^eZ�M�"��ss�&�����l�M�٨����y�ޠ�,N�Qi�[�����l�k����e�Ί]�>�]h��J]l���c���ЩZC�����9c��=2aj��}:�4�:�>�z�abی1�"Q
,��<�hbY�E���hq�yI���g�Fr��Q��D�'�Y����IХ��L�k#�~�f��q��#�"g��lAH����c���p��yչ)��Yer��6ηA����Kd�Z��փ�{�[Op�"C�NĐ=�*�>q�����R��DI���頿�M5N�.4_���J��0x_TCx��'b9�P�br^I��s�$Dx�U0���q�}�f�|�P'#4t����v���/g��n�s5 1O�Enz��V���#)���)Ά)r�����`p�}�uҠh��T�����4���+	<����&��!<�t�o<�ĵh��;_V��h+�` ���ΌR�M݉�Z��"��V>�l/,%TW$��:sb����_,�q���֍�?��h�s���H6�;�Z���J/b�3��2Hs`��]��c^~����rI%*��]c�b|`%�
��x`ó��AG�"m�~�KÛ��ŜJ"B2|��U߉V�J��N�9�ݦjxV.�-w�Loڪ��t�]�dֽ�=	h ��+��$��Ճo�"����=,��%��h�s��&j�&��0�%�:T��,]k���R][���}3oW�2��I��&�T�"ؘ1zFd;�yQ �ג�E|�0.�p�ԄN��4�W���*[�a��$ ��9����*�Qݱ=%W�Xz*Ef|8�uIq2�zDU}�����3����p9Z����or��p���=�˯;`�a����<��Ţ*H6�)�Q7S~|[�#)��C�O/�+�g�p.f	�k*[Z�|c.?�&M=m�:
��G���@V��f|)iie߿++**r��"[��f�}�[���m��߆��^aY�J��V������/ �sc_��Q5c��ޮ������k�ױ����A.#��e���0���?�;ay�5m���V0%%eINTF���M{|���-�R"	�C2U�� 9q��_�Z�HV���v�Ԥ�7݁��Ӈ�\�	�Q-ᦨ ���Et56z�F����OM��742�!H��~�:���0�ʛ���gh����X�/�V:K�]vD�w?|�0iY���1�ws�B�L���c	�1v��b�%!�'��T9gN�!tֺeH�HL���uSr�[�L��	؃���݈<�=N�J ���"Evvvch^u�k)����
���ɂL1����ؠӭ�QWRGC��or랄Ӓl+�p��x
݊�\�m�ٵ_/�toz7R<�Hx!o�Ԃ���-,�7���ᩓ� �=(�d�|ǟ�oaQKM{�n! Snk�3�,.fu�����ew�(Z�����Q�)�pX��Fc���t
����T��kنC�R�#�����wد�;3�-Ԥ�3J��8F���'��)!�.����9�y���Z�d�X�<ǒd��黽�7JFZF�'�~]�}��?x���;�@O��O��bYJ�P��m�����������Q��š��������jj�::Ӝ���++5EDD0[[��x���&���R2j3-Ɇ#ߘds��v����?�}�.7��Sm(�������I�C,V�d��릕�K*�t�;Q����ip��9���ϕF*P5D���u������S��@&�W��ny��UFVV�1���3}�⮮h��6vp�s@X����3d����������$#����&�dpppjn�a=�/�;/"�����&f�����xxL
�ֿv�Kρe���SOP�7��<Q�Ȍ_�k�*���P�Ʃ*
{X|��I�vS�d�!i�ycde�n	>��wt�zd)��Y�)�ZU�����䊗�BxTt�nS�S�ɹ�oׯ_�B"ˌ���=���X;���f bpt�ңrhc��Է��:B��hN��+��L��FD߭���������^��RȾFi�@ޠ��6 ���i\i��,�}���""���<��{&y@&�B{u�2b���}�f��\�$Xt&�#/u��0��Y���Jy;�M��5==��
>yt¿��?s�~������mS�K¨�+_r��ή����֤���^R��\ԫ`§�3��uu�pQ��NR�k��Yd��������U"b���c�?Z`nl����m$��ȇΩ��cR�^�W�>zu ش`��a	��{�;sy����!歁�II��U9ii%}l�f��馊g˃@� #7�-5Ӿ�l��b���n)}u5� }��=�̀@F��ΆA\L�ϳ /ٖXgj�B4��w�H�A�5��zw�����S��֖c�ߕH"LkcR�[PB�		�>u[�sU͖�����;��W�"��~7��ݖ[���H�{a����Ey��xS���1�F�Z195�n���~+�	��[T�Q3��J��cSx�ޭ�>�7svr�ɖJ[b܅TV���n����s����w��j��;�g�1�!2�ul :{�[;gX�-�����)g9%�n<�y��*qR$�xg�#�����"�aճX�j��N2��=�651Q������+� >�m�_9�]��jDD���ܳ��:��[$������%&�GU}���	<5Z<<�$���b� �_׿~���K�nF0�*��#0�2�)�舣�=�lIU�H���ӡ������Jss����S�)��6L���?X뛞�o���X�iB���WjO=����|?O��t���S�����\y`\fc���@����/?�{�𹩩�{�7���6���=##� (�[���������h\��[t�
�b�8i���(腁Jk������s����E^r%��B��O�7
�gn���������LDm��QO&ho\;^O��c�����[-�Y�����YFՌ����D5UU�kǍ�ShV����\`���"Z�%�i|��o� �@���fD�)��\�Y$�Bm�/̵ָ����PYb�Rwɹ��]�j��޴���9oprrJe�A��cW�]���g8'2QF������4 ��2����x�3j�`���3��E���� 4�.�9fd��k[[�Dm߼.Hi�<��Fa:�.�u���h]7�''v?+zP��"��7���JfX��%����;�lnV���|��o��ӱ�l�EH3S�LEt�	�\V���n%�Kz��3�O�FJ����^Td�y0>�PoQ}G���]zZZGo�㋚�8S)�Z���Q3����R=cc��ꛀV�8������T'Ұ�1��W�R�#�R�!��VM���4]����$��S{�G�kS�W��ͤ��N���:%�"�
�������a�t߼�����,n�9�N^�g�ԛ_�H@s3pW$]vI�ޢ�7�'��Y�nv�O��/��k=����.�ږ����ڨA3��)��ת=�s�v܆�V��0�
�=d6/�����395���-�� a��p�� ��9t����|q�Ν��
�8������|��Q���r-�_�uw��Ǧu�w�kؙ\��̨V�Fn%{E�4O��&���p6����9��M��J!�`�;��L�Դy���X��n�ͽ_�W�4�p/2<[�3-
yv����|7H�"p�������Y'#�|Sçk�9Ms����>���[ZT��{��� ������x�(�qi�k�/Oҳ��J]�Ѭ�:NP���|�c�d�oW͐v�"c���WT��}:��������6S#_%y2�����Lz�̌�	 ��s23'���^����~��Ξ�r����9@�ۦO���ő������U�V���|p;�je}�H�>C'�Q�N$��m1Wk�p	�򬾈�t	�̕;Z)�����ǓDT�ػ��bOb+Z����/7Y�|��TZU��P\hm�ņ�M:;��$��2����ͺ����ֹ��'nS�`Pz�Y�s�o�l�^.���J��d0��Ч���ٻ�3w���ڦ��PWw�����V,�6o�xN�o�Ҷ������>��77�jco�U|kuV��c����K�~5Ӑ���i[p���m�xZ,�5��D���?�{��vo#�z�5�=��rOLL���A�.�;:�~���+���M�$�QCs��������#�ۏ<����l��jlm9ﺕ�Zxс���zC�N�)��֙$v H�	��5O_������v�R�9��T搖��q�Ѡ)����&@a�$�G|X�Ŧ&,(�ld��S�����e6hr��MM�C"���gs�� T�����!��Q�@�'�����p�}0�y
���)�T��n�B����� ���pM f�H+NN�BBB�P���v�'����V�����G�("���h!kr�8�]���\hFэ$���������=t��S��>a�з�ml��0Sػ=[�/w�,NF2���K_$�t麅�݁OZ�(��{�"���sNx����SS�@���|��n%޿D
|������q�� �.�^��WA��|ek�*���-w��h�oqE�a|���Dwgg� ,�VPb�SA[[{�h����n�+]I��96b�̞�ܣ�e�M"g�F�3))�g��Q,����[G�o�W�w��%����m]7g����/����S�PH=�
�k�r�L����̅�e�	��IP�����!�	<ʾ�#Yxm�yG�� �p�=D�1t��HM��>ۑJ�YSo�o����I+{� ��f��̻����Yʪ��P�[{Ҹ���3�����nN������ଦ"�_��S�
�a$`��)[� ��d��h�A@&L��K����H��0���� 6Sa�h`ut��Gf1\VH���Ѝ�(��I��N26@n�/��P6T	�h �-�k�L4�n��y1ӌO<h�����P��w�yuuu�V_\\L��& �k��6�����#��4��~ ]�ЙK�*��A��o9�~����Ф�M;Rj����͜��T!�+�[���g��� g���&1o,f�����^D�̌�������J����o��-T��2���>FF���S����RDp?�5"��C���;�d��:Scqo���
d���KT�X�@!���L	���w�/�Pg�^[t�7ng>���Ą΅qЊ�2F�o�wI@a�5�4u�f�ַ~��������	�Ɖ����f�0���X��^J*M���]���^��~���a}z
��)�K�o��?�x�yب~*S������n,C�qa����B]��&6F*EX�|#� �K�LYB^�%jB���}�����3@�24�-.f�M�������:�/��R����`�3B`�%6|��V���}���`@X6�/]?^��3>r���V��o {����:~w���]e��W�5Ǟd�����S���R\�7���{34��͙<�U���Z3n�Gگ�Y��YC����3��	њO,�����[	|���
�ݻO����O����w�*"2���Y�4+�@�H�I�� ��JCU�t�cgM?��64'���d$��t�*;��q[�.��H4���,1��&�Ў�k�Ɖ���p�Z�`d#�K�V��m�X|@5*��2Y��("����y���3�7l�2wW�1������405�Ϭeq���Oލ��5�V�`d����	��nV�Ջ��F��\��ųn�u����uo�}6�ǷWK��r�� ��)
���rX����u[�T�74,Y4�f���1W��e���`�����g��)�6�����fԕ�,n1�_�?��y��\o?��S#"��^���{��B^���N��xI �fe���s۾~�h1'[�]����Pw����Г#�-�(a3?�aD<��X=hP�̚���Ȣ��颍-:W<�~(�/���|V|	�Y X�"�e��9������F��^?�th�Y����f��߾��x���ԡƃ@���[an���a/��e����wl	��c���ɒ�j�.gr|"~g�Nr�y��I�^A�"���(�OR��=�["h=�_Z�}��\eX
�2�� �H��V�,v� n��(D� >كy��
6n� ���+���6�2F,'GG���hkp>�yv�훶Z�o�{��^F��x|z�r��R��1��W�����+�Y	*|~bő��g�?u��zO��.��I�T�&{�@2x�MZ�%�T����j���~GP���j�>>>\�ԣR��O.�SMv�AѨ�����B�pJ{2���C	���v�1��|���Vnyxv�����	V-Ҿ�`Ƃ�.̠���25;z�{h���zu�®�� ĥ�o�Q3�vt��LDD�(=��Ӌ=k��o��Y;8k=8�8
l5���;<:J3W�c��47C�[ZVU�"L�F�5��C�; �K�U|xkHᜤ�4'D��8����+M��69�
��{�c��vp���s��b�^�]X9L��2��D�L�ō��B�;��]�)�a��x���:@�i�<x�̘��)$]brNNN���F�'
�� }�V�γ!��w
 �P���5����۠0Z�n�a�B����-��CC�]�ݧ2�*��8M'wꩌ�>L�]��4�V_ŕ�=/$?�U��9�}��w���Q�/�%`wJ4�M���%;$�[�0"N�G�;�<:"Q
 #W2�.�����7^��jm���2�zگ�L���bN�X�>���ëCv�]���$b��pI�Ü�W}=~e�q.ퟌn[#�=�ˉ��,���/y��-��?
=kG�{y u���d�EW�`�0I����d�v(N58[��]�M�on�3�*��D��3��zk@��|�o$I�N�~ky�s�v~�i�!�S���F=N���Z��	���Sup�N��N���q"]Ȟ�<kyb"��Q�(�~ww�.������^*�,,� �rʬkiM�|f1z���R�v���E�>�w�߄��V��քߴ"6:��K0�{ZZ���x��'ѹ!F���&���v*ï������?�,k�Ov�w�n���a����=�ezPϒ��t��2��f�lS��Ohkk��׷pj+^�u����s��g˗H�`�B��d�P���ڻ{�+����	=��*�l��x���xأI�{�B/ٌ��^������%�w��}��rثg�Y���ۛ���^*�����"����F�,bf�@V�|~�$ku8Egd���R�S��\�[i>���-���F�U�?��)B"� ���g�-^+���������訨u�2K q_`�H��3��z��|�{H���c�%����å�%������ξP�8��~���a�C^�s��E��.�j� �7l��Z��"i�*�s.�C>7��h�m������5�)���ه����p�В�$��� \�39�>�m������t�Y?���b�!ٕCp�j�ʧ߿�%$*���pTQ�؞��P�����ga�G�b�
)))��=q���σCC���@�(�c�h���-,*c�T�SZ�	�����)�e��Y⻿L�؍6��k�}�Y�W ���>,�񨚼�&�qnշYW=�[��g�)��4ۿ֚���j�����}��e��Y�i5��`�[�M����g�WG���>�ճ�]���
椄�'�����
�_��~Vh).^�:}���#��֯�������oa�L����Ɩ�ؼ��u�
�?�g��l�<::��lLOM���;�qjf�nedbB�A���b�,U�
�/|���ʑ��f#>3�xJ�m󽠜]�#�QB�%�
��J-����z���Й�f:Aʻ l��NhZ-ط/��Ϝ.��{(q�z0����S�[h�U�H�5W�ǎ+��T��h����%>;�G��?��/�&+K�����~n���(\�m�� M�^�%&����7/ ݎ���wu�-5�:88��e�=T{~D<��b���9�j�ʵ�8��� ��ڣ�%05�gŖ�m�{�v��gg�LI�1]����������G������싴��<��Ћ������'��?^��m�R=L�))���w?�Gv5��&/D%�	�?��;��둞��2~i���J� td�^��N �/�:'��X�uתu{oB<q�BU�G!)��e���d`0`��x暐pp���q�@iu](�`0�pMӯ��>�)�4�M��������p� ̚}~�u4��
��od`K��1�L��۝�������ǈ���+aw�R��z��΁�վ>[>�����{�z̖!}���9��ᴍR{G6N���E�e�A�\N�-D�p�Ѓ�z���M��[�r���:F66�w�6�� � �h���WHN�d�!���d�0�F;{/
j���_�
�������Ҭ��u�,�`ȴ����;RQ�1�&����N�����v�O��E:��5Pޯ)3��!@"2�������LNYM��)���ޯٴ��j���S)����X k+�7�[��9(I�8��H�6���QA}p�R��eG
�Z�i�%�G�81��:���c��[�n�P8��pi_J8#��h�>J��Y�k
w�dy������e���p`"'�׊����!�du`H[�%l��.�qq�G���Ӯ�:��e~��Šs�D�7ٖd�fB��ˌ�.���}��;��-w$A�̌�lsm̶_�$��{�r�]���@(~���?�gX��.!�7�\�)�>�Z6n���;�?�v�*�E�������#���_��x��U�ܒ~�3vxx�g`PE�o`���ɾ	,�X��$|r+�k�-�.��`�'�i�yW�˭�%M]-a�r1+�u�K��S�cD�.g���5C��Sح?�t٦�b���g˽&gp��]|P�y��������K����N6�^F��ܹF]�0숰�RK����NC�OJ���Ԃ���V͖ML����Z�:p�Hc���"�h�բ
H*��R
����G��vڿYSC�Yˢ(HYk���>���� I��B��j�ڑ�{%�ɫ5_	��C��%��k!�q�̤N�If2�)�G���s��Y�Z�+�q��F�:nZK��z��+�4ǝ���a"��U���ů���xX�<�������]f���P�	�
ُ,�0]�oG��Z�&
��7l.b���n��
?���UC��7^B�	R���?q�]���m�(��Z�@��<���짽�F�f�,hu��C�ķ�E���Vt���?��g��.#�`������J]Ϗ�����jèm�&�M�� �w�3_`���j)I)**����l��W�tu����0?��z8 1;��E4t����m� q&�.@��\X���9:���;dD�J�5�c#�VdT�bƒ���[��F���ݩ+U=�Q�Y�D���{,II�g`�~܂A-T���|���]�y�Ƶ��3��P[�:�CVB�@��<,��+J ��E�U���M�d�g8JzL`�њ�e����K����E�f[�sBa�+Y.���=X��hU]0�|���i�>�S?�i���U��:5�B�y��Ex��0U��C����Oxt��CTD��n��͟t�k�s������}I����Q��<^S���
ޢȟM�X'�O��"�M�Jra���{�l���Z�J^�v��$���*��V�y��鎞�>WNv���~Q4R	��q����|��2tTc����3O�{b~�T0T�6�6�b��d�*:��d��@��`|3��N�����h���xlj�[R��][E�Y'�A�~U�c'1���֤�ƫ�r�{��SO�#ˣ���>ǘ���ͱ�Q��u4����L�vQd;�=���:;&��������3��Ĳ�Х�4�����4���@&o~�PW�8�u��!�D�BKZ��n���N�23�5{�$�u��D�$zڋSV[���k)���	��#��B :�/Y���֐��6�WJJ>��1qq��MM�����n~N4���ˡ�����E� ��q�'w�	3�8xL@	���ܟ=��e(P���#5t�aK�����?J��γ�$���*Ô�G��t&g�	8Ε�;_�B��jl[�a�����Ҭ�P�������dzZZ������,��(D�n��Ĥ��1�1-&(�O�^�X�hj��@ܼ�N�w�;@[eA���o�)�(Ұ�%I	-�0�W���%0)�0	j}Ǐ��u����������w��=�L�C���:9��ܣ�&WWףX,Ƿ�?*<),".�����v����(@	�ȭy��m����ծ�@���
�	*�Oe:|7?Mh3�����-���D�k�e���0��� 	}L� �҆0�1��-UW~+PYAI��3�� r�Ц&� 7_�g6 �ه_���l �HlSss���?YDMKOo�D�H�d���f�ʯ{� ����f$R$J���>�=��mA��f��,��]0L�閞�B���x�O�wSS�G�w�L{\�H0S����&�����-	��C4���	����w�{�,�������3���w �E~��O�i+..~� �<�R�6��Ի��g!#I)�U=�§�8��d��(~���M�l���(���΁��٦t)��d���<��J++g �Й�.	kd��{�컫���08���#+�LGG��6��2���a0}�18���Ζ�ُr�ա���m�c'�Κ�Қ�E�j�I��6��j}��ݏ���:���!W�v�_!r+�b�d�VYm�aBw{�@���_W�;l�T���|v�(���.��{ tW�/%Ԏ�"r[[�u$�ȼk���-SJ�Kw��$f(�ٽL�� �֠�|���7ܮ�羊i��ѻ�=wfCV�8D�PN
�q���ŷ��~��^\\ж�4�lo���&122ޥ�ξD��
�,��S�0a�u��# =YZV�V�G<2�=���٩ר
�uxQ�ydU�D�+,~w����!�/F���z���0�UøQJuu'<9�/Bq{R��gmG����j���/Ku{|�+����e������\
�eq6��q̻�~����2TC;Tkk<����������+W?Ͽ�_<;�H�չ����*��>2.!��~��-�'�p�\\:fI���><m!��'qj@�<Z�p�&>�EJA'.{���-Y�[�	ml��d���&� �4rh��������)�m�WtVa#����P	�;�KO�·5�����
�)W�ɩ��#a��s�P�kY]�nEEfs3ޮ�)��yV	I�}�~8;g٦&��/_.�0�J�Ql��	'�+�0t����$����c�śE���:����
;|ph��6�[��FJII������A�ǎ"�(33�$���5�MVB�I�=�5�w���H.��H�ݣs#|��6W���T�$�k(p%�Q(^#�}B���p+��]!xo�{��1$<E���e��R������ �2�uo�}�7��w�"m�9O6�X����kp���M��#�14��ea�S;>f����p�?�ݳ>3{{siB=.�F����i�ꚸQ��"ȣ�HW��{U���{HGP�(R�!�B%@@�މ�Ф%@B�Kx����Ϸn��]������3�g�7{f��W�m�N�G�^�>��0�2C����,		�A������~t�^�
�I%'��a�E���e�>ڿ��� Ej�������̀f��y��d��-�<;����Xe��R��z�M�LyE���YAB`����'$$�#�חu�o6y�V�txL��뛲^�߲��W$�<������կ ��h�-?��x��4_x� ��*��wN�d{��Իǀ[fyhV��eu{��8L����l����z�Y�����I����l�g��cSOU��*Ʋ0�-G�Yd"�ϒnm�Y�j� R���Ҷ��3�b�s �Zƍ�-Ve
�?£M���۷I~rE���j(�#w�3�2cA L������#C	?��t���w�ja���snj2�K�K���F��ӛ-Ɖ�%z�>�뜊^�|$'����$�hy�hc�p����+��C��oFQ���t�)��u�}�ǉm��OY��}O���"�* ��z�eI��|����ȳȚs��A�-�?�e��G��X9:�ʨh�!��Z�V�tbς�F�#��
�}�ft�׽�l��㢝�R���D���g����V����b/Ox �i@Z,R���
�8�^$��e0��VG��۫�Τ�5�ȡq�?Ϸ���� �&����5��u��E��	�'R3���'C�b9v��ēn�+Ǭ8͈/K��,��Sr�و�A�Y��6ķ�Ɔ���e�OJ�
_�J�S��S(���[Vx�꽞�G�!�p�;�v����Qtmm��Oٕt�+������!X ��þ�k)���/��5�?I�&�7�U���	0�3W��w�>��^��d0>�'�t=�3����m�����R�n���=n	�Z�׮�_	�7cq��H�4�5^��A��V�7w%�->���E	<|Ϟ@���|�|	����sm���[����{��&p�]x�sk�L���Ɨ�#�s,�I#k�D��m�����ֳ�_���l"E��討���u.*��? Z���I!����U�0��2Y�y��`�>@�3Ic�*��AO'J�d���}J\+��BE �Ҿ��E)��j8t��;��ƈ;6Wq�,�<>��J��|f|[1�����'ol3��׵�g���D���[��CD<�ޟEſ=a�UDY���Ŀ��݁h����ٸ���vZ�ś&}m�=����e�0W�6r��R�����[�|��B6�9����ƛ��K�[��G�5��_����)e9�g10�D��[�D�P����Z���j�Ъ�j�5���+�)��\|:�P0�}��lH�� U��bk��%&��'��)qޣ:�G����Y�HO�'��O퍌�I6`�S���i����'�ݬe��������`2P?��A�<�>1���%��Lw�r���qD�\�a��bA�y�y�'�������o�r��I��qjU � ī>��#�(Eo1��d�C���*_|��6;�z�<���`�ˮg��U(M��{Ǻ@I���S�}����Բ"놨���݉	C�{7x��i�O�AC�3����|1	�H5'�y��Lf����>�ax�ue��D���p�h���)��o�߰��5�ZZ��9)����(b���4�� ��_�j��'C/y���{j4��o[���+F��G��U�A�&�h�ݠ~k�g9͝��~!/kr�o��#�It��\㟺���D��Ԣ��"���d�R�(�w�&�0��C7vǙ� T���'��]0\�}b����Z4MA�G�k@���[��(��ыQ���*L��$�$c�f�9�d�}jt�ć#T[w�ؕ�rDc�K�e,Bx��f�A�P���mJ��G!�����-~�l�\���'�}[#������[�!Iov�@ēl���Uq�g���^$!h3o��7'Nh��;�1e��	�jC�6����n�h;��T�0�%�h7�/ ������/"a���♏[�T��
|W^��Y�j0I�]�T�9�0���(<'Rc&���5�<?t�Ab/̆<Pô�֯K0e_��V�������k����A���q��>nƤc�\����T�:֕#%�Ԙm�s�����G���]2I��� �R�t)�Q0���bk@�0��;s<��/�E� I�,�*��'%۫]�'�hhn)(ĕ��w��^��������L'�#g��fF����^������ظ���o,do1�����(h���M��3�s��oB��M���zƽ�w�T]���K��ܫ�SwF
���E
�ŊQ�FR�K�6K�Mzr+_8R�{[�$X>��%�]�c���<6
��۠��|�l�HbL��d��Jۖ	.b�IH^l��kj��q�G4��3%���)���"kV�,�gIr�.����>XF�愹�({���c�Х�W�[]�5�C��Z����I���_~_XWx�R���:W��2p)��������x����^�k��Z�1*\����I5d(g}������:N~�<�/4��Q�3�+'�P'��	(�/�.����G;=g;3�FԎE�i���a!qUaR���
Y3|�͜X��^�>I���8jq��BCᆔ�ZX��	��(k�k�a�g�<���fW��%ÏTR�77?�+v�	4O���GЃAY�y�����w�Z����O����[��#��Fj�sB�w'����]dTh,��4�x���������#�	9hn��7�?�����	� ���"ړ>#W�l�}15��ͯ����6�mQ]����&�:Ȉf�N�Io� P�[��Fa�ѡ�;�.�)u�@��U���=��6хt� X�Y}��Ȥ�HE]D�Q��"�¤'o�#h�&���V~�������[Wƥ��t�8&�&��U-���u52{V�Y0�7L�Wt~%���^C~#�?��Ʉ��DIp���W4zm��=���4��:�	�(�E�~R�ৣ��B��p4��i{8�%�*R3欳�=���>�Fl|�t�*Y,U���Q���4�)�>嵏�D������	KD��f�r� �]��_�Y��SsRS�1j����8<Ύ���z�7Kה<��:�����'\{�w�j�X]����பb�$����z�3L�@	����6w<��o"`u�TyM��1q�!g>?�f�[�;��������X�Q��m@6ih\.D��E���� �_j�`���3�x�����x-���^�;���������)�������O'y�Nt�Bܱ)vk�8X[�Deo�����{QxW$��Q6S���t\���`���+~ת��ᄬ&�����p�^�I��Ǚ�k��o\Db�8
.T1C�܂�t�N���rF��($^�a˵'i��b��=2�cc(R���;�Ɩ��>�?U��z�G�&�+OJ�ZT�M��Ϥ�Ѫ�G���W�oU���G�N(�{�vHy�b
 ��ڜ����Ь{M�;�W��'bV�[����U�Hb�$Fd��h����6�Y����;��ibF��E�p��B��Kv��)ׁ<���$���B��ŧQ..C����O���w���z�V��d�+J]	�Ǘ�b��(�\಻��4Wq��WUHGǸK!���g~zLژ��K��ݘ��`f~bD�jĶo}�x�S�~��}���z���#�'�����hF���믭Ѝ"�E<�#� /���<x�4�A?�u��m�6*eQ�k)��쓌�6n�f��"W�Cé�Z�`��sI���jHd�DFB%w�����'���5�ޏ�h�r�W���hjϱ�N*@�&k4G�L\��aL-��||��BE4.�,�#�$�;�����a*��X�kT K��2O3y,Vc��z�`�L�`l�[��8?H^�
�ܩ<�h(���"{B&H5S�ϡ��ڳ>��=o4[N/��s���L�3�� �D_^�]='�\
q҃�О8�kuN��Vx�eL�jE��&n�D�;�����ٶ�=X4z1��>��m���G��=��뗑�=�,Qa������������:���<&F��%B�Z/Z�(����/�\0��ss_�=î`�z�����fIJ��+�&�'��e�X�i.*�'ܐ���+�8�>�}"Lv���ޕQ������M��������?�ݩ`k��]_r��*~�����HIB���==�v�\�U�Ӛ�/���C/�+�������م!���yN��Q��3�ȿ��a����/o�ȺnI��A�]<�
�b���,�oT{��f�o������d����4�w�?
�5��H&��"(A?��=�`
������|{�jc�=��-5����s�7%)I*���Υ�d���ڻ�N�ͨ-�'� J�(M��W)��E���|�!|�#�k�%�_�=֐v��mn����S�׹x���(����w˜�i �rS�L���Ј|�N��Mq
�[��~�.�@V�j�#�Z�Uzm���)����o���������I�s3������W�����M�&�2<2�Y[���{�-^G��E�*%W������A/|�Q�|/B���F���,M�C��DH��Wn����'O�l0�-����cm����� "�%��}����h����ml���t�9��:C���a�f;�|K�������峳r��O�L�|�ud�i�&]�'V���c���Q��ƾ�ic��ʼw̛o �&L��)�Xt�,����4�B���ӶY��k����%/ VѤ�M��h�Izv�-�1�9���D`��)��)�L��I,J�4 ���η��X-i �>��T���昌4�N�`��� N��#-e�Ŭ�}�p?�Ap�f��W}��A�O�"�Y9K�>��5��>=�����c/�Q}?;�~k�z�9�nf7(�,�8�tv�C�P��`�5%1�RD�?uؗ�O��g��G��z�r�D���5T�)��6�#�b]�V	�m�4�fgk��?�~@lF�c&�i)U�A�#u �js74'V�����-���j}Z�$8��Rkd868�jI��a�zh��&�_*'l�B	�����a��c��l��8��Hu�|ս�S��?Gި�v��fJ��x�=��\�a٠UMy��0����8J�m�4�u�����az���dKhHž5!�d���V�e����t�����H�Ђ�Rw�wc�`a��A��(\oc���"���{���Y��X����F��n�2��!M��Y��K�Ǎ�N�5�0O2"��
ߖ)�������׊a���X@�pviBy+|a��%�o	�|����g�R%�mn�����)�x�U�V�'���A'0�|#V�;hN�-t��	&
5����-7xM� ���\�`�`0�A��%���u�sP^JBW�*��w����&�`0.���vz�$%Mz�o~�}З.�'wc����y%ó�4(�
����6h�9C�>�Q�0�����d�s�����y��!K�
�c�D��y�a!����kZ����O*Xᘟ'!�P��]����vPsнqeO����_B�Du�)���a~&iÑ�o�p궕���=�r���K�5,,p�g.l���w�[|��Ò���HF<!�т��?6ϰ��T��i��~�w,������Ɯ;�_�a�'��B(�ƺ䐦볖��m�\n8��o#eu�I�@�ι��ҵ�T ��v_(%���)�:��ٚu��G#8���y�}�D%��ƚ���ޚ���5=cY��&�of���'Ak�g\�u|xk��KM�ŋ�7�ۯ�C�������x�Q&�lA����n)�UQʷ�F�ˬ=2m��Y���e��1�E��S����u*�f��n�=�a�cK�V�N"6F���g#&�Y.��/�K�=�m�۾|F���Y,I�6�Gy����,�1��,bZ��A�d�dOV�m�RawΊe��_s�t�gL��V��>�A\_G��^abd��נ3��mG��ޯ�73�웥�(}�Jڝ�t8��.���!#���nG��W��esf��߻r@��*���E����s�j�����h����^�[L����P��,7g�D�4%=�w�{�����&b�{"X+ ���(K!GCP<���eRۅlM�"ϒ��l,�>��T�[,��?^H�r����\�/�����E)�o�z���x�ν�*��:@�湦�˽~��׿ 
2E�36�n�,0ȂӞ�sc���B&[�gI��SN����P`�GVc��]��S��i���>��Vbh�����z� ���@��M/�6��y'�8޾{/��fk�A͍��g&�V����=�n�Ȏ�q������7~�����ҹq��N������G�
�a�f&�Ĺ)�d�da??l�u-.u���� �����3-2��F�}�Cm� A��.��P\��3�Z/s�8?m��o�ZHgwq��l_<���-������/���SA6�;����+��sl댏��4|�=5`�5�|b�����*S�_��KH�"\%�bX>��F7z�0Uf��?aCl�mIeN�d�����!����3�e����O��ۧ��+���VΕ�ۄ/���8D��6� xK��i�T���H��,53ʈD�<�n�&���Y{��)�|��s%H��!�rdyEr����`�ξ��h�~J�H7N�7�x�K�Drd�aR<2	��a�����u����bw=?`�V�e���k�-}����JӋ��f�����[�9���L�<�΁�������+��v�U�b@��� ���`�ca���=�2/�0!U9��hn�q��+8�0��Z�Ø��k�d(���p��V��M���u-�͵��2~�g�>q�l����_g���y�Дұ%6�W}+����5��i����_܄�gc8նd��\.�@��y�3'�1O����ONa4g�哦���t-�X�I�n��+��!	���-�#�晋�$޴��P�����`��L�����XG�'�DEz8��śE��j���!뵀A]o]Q�?�s����<���+ϖ�i���PFm������eb.e��Fn�A���sm\ޥ���x�9pw�a�G�kG�LVp��2�����I栉���R!M]J��_+n�Au�� )RG�L󓂑K�*�n��9�l�'KUg#���GXH��ft%���U(G������ڗ��w�ql��D�udx��׻�e-+]p�2�R���Z,�7�j]}7�]�i|D��+�A��ZH��)X�R �e�R2����إ���G�u��ӑt���T'���Aa}n���	5�4�UZ�Q⬎u��m��RO�{wc?����ب(x���f��l+��/-��z8�02��I]�]��{+Ti�8�W�	6�<5�У����R���"T�Ү����L��a�P�^z����(�Ѫ���|�{W�;�i�S �\��_���F� �&e�aڟ��fA,0�焎$��r�5���$��"d����U&TG}��������l&��HG[�_W�7�I�|�"�6�&oc�������͏Ń(ƥ�ä}�_�n�����yF3%w?A�q���+y�>�m_г�D���UW?��V�V�V�����j^]��w$O����IO��7Ä�Ǐ�3�ZZ#o�r#�tZ�@�e M�M6:��!�Q��J
�K^���݄���J ve|�3]�
�_=R������1���$Q��c;���~mLԑ�s1��chx�>ieӵ��>�W^P��G����:����xpTq�a�[~�����>z��sc":�*�8~���fQ,�Q��ه�D�?��/�U�u�DiJ(^.�+�ikY
�j��Үr�_�ǲ�\e����f=�D��ѯ)�Mb��Í�쫀�k��K�+[-cw�u�J2��#<÷.�7L��'�8,_������z��I���s4L�	ڈ_�YQ����}��2R�iM�J�[����c�I��=q�v�r<^9P��5jsѩX�������AݚK�!(�)��i����A�g�;|�����4__��|�]C��v>O��'�>V�S�wS����,��&���N��?(§�>F*�&��lD���Վ�ܕ��7�G���lO�K
I��w.���$�PO
��y¾�G�r.6�9�9���W��%�*�}�.1�
��ݴ��#�8�P�4�:�,�(�r����̓�t�LU�2H�?t+�mNN�0Q��
�BP�R��M����'_P�l}��4��e֙��O�4W]����"�ErǾ/���n �Jx�U�:=!O%��˂.~GD��۰m�D�{�&G�J%�:LSQ|խ���H�o��r��ݳ7=YgT����=�o�SV�Y�U+��A_��I�@XĢ2��J@�����r	�2�Epײɟ�(����g�m��S�%#�Ǫ�Z����
<�vO�y��;�&�(a����c�{S�h��,/%\�w�T�Y�r%�i�_l6����D���#�4(8��h�t��I3�mzd�D+�$~���әW�W�4`��_�T.Q"�T��b�� ��N�x�\i>�Y�-�P�{\�U�닉ŧ�����_��=6�>��n,z3'���W::)T��U&N���zCoҭ,>��+;����ėx[��fd�c�O$�C�DarSy3��g���t�+-�}9V!8�y�h�i�'x�8�&	#�{�hD�����P��xsoh\��/��#�]��=�%��W]���"���I�3=�Ap��i��>�_<�_�"M�J���S[���P���985���b�r���/ȷ{~__�<|�����i���͙L��'<��A���,O=8�Y�����#WA��	֡��
q �+�}�W�]8F�����`�`���pJ�:$�!4��Y�F��#��'�F)��<Q u�����^�M �M��ր�(�s�t#����z����*L�����о��h�#���"k)�77d}=d���P�T�8�0����b��P��oO���� !��9��%�W'=�s���0��s3�%�芔�O��a+��*��ט�Wv����3��玡1��Uk�n!���H^~�"6`y7���1��AҦ���3B!���2s'6�gҠzmu�gt&�K����6��`Ps@:ݷ��M�2I�r�mԚ�L�-X�P���?�zo=u���2�=��%͢ga�k��+����S��)(A��O�.�^)��E�@�2ψ���DmX �� ����ɚ��LZr���C�G�[B�;��	7�)]7�/<n��	@�����3�(�;c%�4͓k#��^���#{O�WŚRH�R�^�s�=8����g8��\d�$m��o�M��Y��dR�Ϲuv�ʾ��5��Mp��Kx��AR��k�*V�uAs�Ci��_�+F�i�N���Y*<G:�'�����
7S��>�p�5�Iޗ��D3G�TҎ���T���	l�V��������?E��Ф�&��z�|�8vNe�ۭ�X `Q�z�<Rj<���=�	"q9��9Zo��2� �E^���>T���۔�h_��=�g��\'C�  Q�hM����?罋� 	o̇RkYf���Ŋ-����A4��Y��d���&��f=���&����Qũ�,cQ�iaJmE�O�\&�ǣ3�f/�^+7�O[|���5=wg�~��<�w���qF��Ҕ���!�%�k����r�m��4�����@15�� ��Z<�Aҏ��иo���W���yXD�'.���(�=���/��-rwrh�xr�1C��Ay&�}z�Y�jV�>�8�ڌ?'k�G�i)Y(�`� 2���o�|j֟.�W�X�vp����N:�e��]���_�&>�B���K�~u��+�$XZ����ܠ|��㗛��6�m�X߿{��ӺX%B��B�����Ӌl�4ӄ�e��Y���Of�uz�m&��UV-9��L<��9_׳�%;��������� �0�|:뫬���ZW�_躀ʸ�!8�=F�]���Z|^�������RLe�&�(R�,�Hte�g�WC�/vT��Ax�ԨΦY�dI*"�E!��K�>U�fM+���pߩ��j�r�1b ��񶫹Y� �G;�r��+] =PÙ(B���9��_L�$���tQ�yֻ���d\�����m��J�ӊ`�x@#E�v�fAv��v�#m]��2������\��'nX�)��x�z�� K����y�6g=�"�It�.�ܢ*�𔷎@�9���ao�h�j��'��4L�
��nAɥ��SQ�<Q������̛�f�f����	Q��+$���j�\2��=�����mU{ho\�ܪ���i��i��PbyJ{������aG��.&���nS��J+�B�ED;8#�Pv��DH��l7)�\��m��f8�%�
(h�2r�����K:�F���_F���b��46�W��R&.=�1cb1�W}.����8����4�ӍV&�0��\����;jJ�6�66V�8G�_\�^���)q�xh9��[� ���1���W�4��Z�QU�oy��8��A`�����H-�����Q������%�F)zE.�6{�����3SZ>�Ҫ���`
�:O�d@�|����-yVI�KN
I�r)��	�sR^S߭��t�2&j� _h89\��~�%�!ԗɌ��(V1�,=`�&�mپ�[���\J�6�:y�Ze��[�����ڛRn�,v�oʎ�\]e�-�	1�4��/������=z��E��0\��"y^��$�
��v��b3����X�m	���]�� �"cN7y�����qJ��ذ����ъ$T#��"^�۫�V~���5����U�,����?�a>4���z��#�I���U� )�+48�E=1Bp�Ӫv��"kIIv�Sn��s�O1�:��@��i�Ok�̛�~*��G�u�W���9g=���������ζ=� i.[g��N����d��h��'����cm��8��X�϶͢+��)xɳ�œ���]����l�%�mκ�h�^�|�ULTDgNk��/��D��q��	�孤K��|�}ԁ`>6�J��9�5�-T3���P�ؤ&Dc������7hβ
~ߙ��O^w�Bw��ۅ�F�L$���G"@��������וT�Iu�籷�1�V,�8�-��`�^G����WL}^~6��X,�Ӟ�0��av�䈔dyL��[	�����r�]���kE�7�d$dPN,��F�;0�΄�)�}\�q��Ky-b3�L� iA \b�Mjo<2�����0�mS�b4�>!=ݓ%����7^�-J�lrс4=n���L�"�<����W��hʉoL�Z�k�d#���_��A�=��y���52:�)JAs�E��z�<ܒ���ڌ�$\e��(�7�̷L>l0�7k�!"�7�F{M�dsmt
}��(�z͘���2��P`;�adn����}>�f�⚲g��$���Gz����r��b�҇&��"�N��f�ٸ?��x6��آ�:Fo����\�X���rx��,�k��2���2knh���g��K��y���u�{��7̵٨�y���N�_A�Gc���{�o�7�Њ�)T+,���G�4���(��j �w��+�y;A_.^�W�(P�t"� '�T�.��wT]ƪ �4.�f!�G��M����Z�m�_��'�}<;�ǂ�Ժy�g;)�\��zt�uYA'��΃��k�D�'7��'���FU/eGE��$p�H秥��ѠM�n\�_Bb 7}g��f��\it?G�<�?-��c��/U�>U Ӂ����D���8��EUS{;������M^�X�v{�J�`� ��&���>�"���S;OX5�e�x�u��d����V\h����5�=`V���r�i�G��~-�U��%����1�eņٿ�Z�_%&���7+Z?��uWm��,V�}�F��NR:
lZ���P�5��R^�c-u/w03�N��in��y;JJ��)do>q%_��e�м\��z/Tg���xa�|x~��;$�"K��%��B�n.��DRPXcl�69vY�j+&����ru��v.n�&���QD���Ye�11ü=~��;���N[�W���h<�x�� �w^ �@�έl$��}�iT���)��-V�Q�{Ь'�*���Zk\�^��ִ,v�W��{���åb�r���sU��aq���J��y7ҢLX�K����f�ZWʗs�ck+��Λ�4��':���x�2�.�:k�f�ͷ��c�*�T��D�<״z�m����$�*��Ơ�X��Sӓ�˗ E�(����`"������8�F����/�W��O�T(r�������(�x|h~�Ry��CZ;��-�~�hP���$�h���U�U��<���s�c[�.1�W��8O#���L��W���eM��<K���6v�,���k��|⁺S�0�E��Ŀ�s��-�
��sx�,i�H���J���N��	�#�8
�-���:Q�-;b@5fA����3�����P��縲}���-#p)�@�[VQ��g3����_���}�2�
�z�y�,�UY`c�h�hŉ���Xј��_��������%<K��C��`�S�h	�-w�q�s^�:�YZ�&�3Q��+F_�?8�l���!��ѫלڹ��>_x�v*�9��G�g7��K�p������h��YS����pq�{�JE���Zl���ꃪ,"�Җl�w�rݼ�?fIF7lUn�a��5�ȕ��K��^B.�)e=��7#�H�J��-�
뭢I�����5(g&�r�w�O�,5z>�~q)Ƽk3�#X���y�~MY����v�~�P�E��Os˓˲��gm�y~�?��&��%8�M-�+�?>XF7<v��1_fqS�Iz O��gw�e�Ie�^j��o|�Nt�ξ�oB
)�5u��7S� Bdd����#�W#���T�q�e��HX��þ3�Z��>bb3M���l��$�bQ����n!V )��z1�D"!��/+)"�mG�
,�g6=&����n������Q���]sU���tZ�K/._�%�(���� �@��|�:�	'Au�g%��.���F%�f���W�?����r��˛��0���J���m���oP�E&�Mo;6XX��@��,��*��[�y*���L�,r�n$�EO�:DOzf��B^yPG��zkB��[��/��}TI�y��N�?��0E � *�#��c+���G^��$�{jZ$��d!h��%�۾e���M�5��J��gxdo��g�����e�{ҽ)�̊*���a��\���j�
5��\� ���P�ל1=�R<) �3�륗�=E4�5��7�!m#��V��H3\�L���Ԏ�:��_<���JjbQ<��>��Kp[���_+嚳eQL��o�AO�,_\�+��hh�_PJλX�)=~�=;�R3���`���s)�薇�!g��^6_��ꪚ y�?hK�Г�؞U��YW����:C`7zr,/�r�s�������Vf��$���_����q�p�I�r-A	��ƙJ���R%c�c�yV�eg�5H�j<��kK*����Z��1�i������^�R�{��dJ&�,O��B�c��Ǉr�+�e�e[/��_�	M2�n����~����T����w����%o�s%Kʼ~�T@N��No�φ��v��z@~�we���9���}�4��{�kl�_�]�+�e�����ͿIM������0V�&��������𵟌�A�~��S�D㬍��^�7��2%?6�a�uu�}��wnvZ��?g�@*��ƃc>r��=6q��p�.�a�y�3$�j�+U���	@fb\K��d+�7S��S$&5\������y �u���� �<�M='Wծ>���ݦ��~߽��q���9������;����H��f]��M1���.CA�L/�m���>�����vc}�w#�hn�H���v$$�E�� ��Wg�n�k����=�O,���OH�Tz�W<��U�e��d��SRk��fL!s���Ob�&���Lk��K{|�K��{���`��%�$�C�������f��/�F����� j�nRw��t>�9^~�R[n�fFE���i<�77:KZퟎ�ݦ��b\�l�`t���pvL�K[#���e�������ˀf4�ŭRr�I{7p1��0xd�>��z��ۙmh��~��Th,:�V�7Fwf�m�$[�ΎT�p�A:�f���������������^��4r��v��~�q��_;��@��~��������Ӱ�+��u���{���!��!��T��<�|��<H��!I�1X��%|���F�C���6B7�C�rG 7G��ֶ��~����y�2��<8���Jn�V�y$V��<.� H�O:O��4��m��Y����(�q�|J�����z��^��c3uw膡.�H�F�e}�Z��׌�騧�����e��䊧�_�V�����Z��ɂBM3s�9�5��yv���f�I�,��mk���g��,=F��#�<5���3�V�䲮A!�t</*#|4!AG��Zz�S �{B��1���t�_�N�z�$��\�I��Έ��Hw8^�r�R�Fug�M�&tYn��<;ۊ,�>��z&kN��ZG�KܤW��3���t�3g��?�G�<*�'$��]���e��t!�z\vs����B��m�@����هټ$ݻ鐶���w{�*ݰ$�u{z�]�x5A�
	��ڜ`]�F��3���*��̟*ۗ�F�
 �'�Jo<��_;��Õݤ�k�K>������� ^C���H����?[��+�x��
��V���Ǿz��������u�p�佫����X��hC5K�/��Zf�`p�]�?SAҷ�H����R�[��"`��_�FՌ��ו����$A�����%���h	p�����%�6l?}���ο��\4a+�b�㰒Z�<<�'�	����O��z���K�1�a@�]y�ԅi�{ޝ��t�,63]s���rxJ�V�䴼*o2��Q���"��{�=�V�"-����V�e�3�{"1�ہ'F�Y2t}���s!g�Xm�*m�$�(��*�k���i��/;h��?�i�i�Q�U�5�o��O䬇&�.'y��I�6�y�ٸ��Ug�6nP}p�W{���-s�n�䔾-��Q ���=��$&>��#�k�����{���dݜ#�����/+|_l�ǷKR�MJX�Ahu���N�[?���!�_���b:W��Bw�5���o��(��}*���%^���V�j#�/�˿�Wq-_h�n�W[���"�n���q7��>qN�׉��P"^�DF����?DI�"�u���������R��	d���VF��>�I!f����������ÖCR[�+2æs֊�d����Kp�c;�td������QJj��r/��;�ȓ 7&rN�?��~X5'mBF�s��e�=��͜����{������iH���q��װ�D�RW�~^����� PK   �\X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   �\X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   �\X�����  �  /   images/edbb92c6-3c2c-4408-8481-9459a63b273a.png��PNG

   IHDR   �  {   ���  hPLTE��� ~�   [���� v� vѰ����� ~�q��z�������h��&&&��mf�X�"�ۚ��$?e�_������쵵����)H`�999��� @y�vtu &n�hhh���b`^p�  8Bn5Z|Ά�� S�:b������B��;6/ >r..1UUV\Z7��fR�/1��bmmF j��L����=��  AAA���ztm������ sט��G� (C���~��|�� .Z I~%  3{����]u�|noR{��}v?{�nu�  (P��  ���{|NV� 5rV�H�Jw�y��*_� 2iy�������� 0u���Di����q��`�� b�5Ol�=�  9IDATx��C�Ɩ�-�z����% @LL %"�#&���( l���6��u��&m��m������5#K��X
��iK%�f��̙3G��T*���V��ܹ��>�Lo퉎�O���5������ F�t�K�Q������D3���1!��ya�k���| ���R��Pl��;9@�"[9PĴ�|�1Z���9�F
1s�đ��!�T�(�fL1��b-c������L2���j21��k)!E�ZP�gJq'!E��3)E�ZR���lþ�ٺ�d��(>�3ׂb�ZP,^����Qd�EAQPEA�1Q$})(
����HJ��SчE��3��E��(ʇE�����H�N ۑƤَ�^���	)��2	O�@9�E�޳�((�1Ţ'{3gff�}��`1[��4�r��T��.g=�#��\.3��f��ق���<���G����(�+�����9P|��v˯S�R�
E�iE&_���o����,�D)���
<,K�H�
��dJ�4��R Ak���=�'��i����U�_ R7œ��c�b�yW�G⃓ͧ�W� n;S�W���P ��:�e��	(�BkyO2+b��1����u\��C5LQݽ7�4�@)$9:���}��}��{K��@���+�S���P|�F�n����������F@�g�{�g���<#�'߹g�n�\��,��h��b�] ��	��8��9�����]�}�S��m�z@�Fم?Cu�LnheJ��#�����Pl�H���B@�� ���[�k#;^�#nG�B�$�С/O<�b��O(����a]�5����t�Ga�����V�G6�Qd(����u"pU�����}��GL>��SǷ4#�	�[����،qZH�ܞ�ዓr��C��ۊy5P���٩�u��;�������yl?"����k�|紑g'�>D/RE7�7�5�~��l~x?B�T4����^�G�_���h���t�����) �Ǔ��<s}'B�3�?y�厡�w�r�"���vD���DՋ��ʄ�˵C�7K,%��(&"EA1J�l1I
�
Ff5aA�@1�k����mڶ}(���P��QR��J"/��BRu��|�'�9��;=U��S�1r����(��r���Y&�)$!��%[7�0�6�tЍ��$ȈI/#�|�ϐ	�S�_i4=�P dڝ�{�B�ޖL�sч�0l��NYr�"@�I���t,`۬�:��l@	J.��r(f������R�նuKL�c�=����t���w`�M��E�	:dEWlk����[R8�%˶��+4�����z�)Hx)P]@�"UK}d�Ԯ���]�(�XV{��UtP?с�+&��/U$ɀ�䒎d�,B�Ӆ��	 d���K����P,/��:�Y��*�w��M�%eK��:�V��}l�@���Nc��
�$�Ćș%A���N*R�z� <	�S�V����T�薥WA�:ԶvF(�Nx[�8��]��Zz�QBa�o���J_����A��m��׈,�u����M�t(�B��D���z��Q�Q;��ۭ���K!�KH�(dP ��i�����A��V!@�ϥ��JɱRA.�� �\&ԧ�D"W�NP#AK�j���(d�B�,i�Bu�P������RW�6Tru!��cƲՁ��R�D��Q�GZ�N(ڔ�ܡ�`lw���6-Y�ڱ����V�ևu�ڢ�m�y�h��W�����R��x�~���(U�ϽmAK���J߀\Q�C�y�l+�ݗ�3��
V����B� �q��&\���G׈�g�P�a�*��zX"=��yb�+�n29�X&[�
u���p ˎ�E�H�����P)�C��N�=�0#|�Þ�}�v$>���A�"�а�m�.VYA�)�L�L;hk��Թ��)P�{a�ȧ��31�B�q)�(֧=���ٔ�0��P4��uO6RQ�]���S"(�$N1|����(�R����Ť)f�`v��7�L\G1�ֈ��_�̝��3w��З��
P��r,6�K%��Ƕ�O�������_���	}gr
>ӟ�Ó?q���L��)x]�P��A��`��((
�O�����=�g��k�<Q)k!��,�6G��$���L��Fuq��C���Ĥ4B))("�$ E���~t��h0=�!n��97G9O!�Rp���(��8�r��p
a\
/�#�.��RQD>	P��'��.�(��������䘧���O�Sl���ؘ�$���-_�8�����q�fp-�`(p\�p
�>�j�)�Cpx�u�\�f�cA�yB��Ф&���ؑ���IAQP|X|{2��M"m��2��n���*o8��8����������Q}g�݆�o6Qi6�n�v6Ѝ;�F�Eoġ.h�>}@�qi_;���	h#��u)C�W?�۳�����"�ۃ�ϐ�����M)hx�R�m�/�#�L��V��Zjׂ���)ƀ�� ?�X�X�c��A�31
Ch4�kq�1�n�ۍ��M���G��]���~��QM�B[S˧ڤu�ͧ���&�a,��[��JA.<? _R�uB��Sz�E)\�˼)��.�B�u�=h]�Jqc������t.^��9]ȗ�F�V{~puU;m�葟Yɘ�E/���/_������zY��XMdM�p�j�˾Z�r�WD�7����.j��Z��S���^8�,47�����Z٘(�~�svR8[W/Wv������ԛO��+K]��x33GӮ&�f�֖۸�� 
�����7�"����D�+//O[��k��b��ljj��à{ǀ|����i��coz�B�����f$ħ��b���R���*ǖz床�@L�ɇ�����˩��Dij�5���W��ܧKAx��'H^v��b��Ś�b���y�C�-��I͋b�^s�i#�˼(�?��m*p[��Ӛ��P��.���~�΃ ���Hh c�y�t2yP@hqzy��w���*ŀ~�:;��P,\���I��F���5���|z��谮���qt�9�G3˿ݸ���c�`��A�������c-*c^��f�	<_�SR�q'�`j�7��+��8�<(h���/^����/��aAH�/��YO�+<!³ٍ�e�aTZ�5����%���+��ΥGO#��E�  'H�.jW����A����������|��B-�q�p҂3��W��@��`�ͥFb)�u&A������8��W��?")2���:�%�.6�f�~۝A�Y�_;���ͺ�K�4�x��ȋ�A�crƬX�p�ͼ�hj���`��T�����OO�x��Gj��}�I-�_�Ee�jW��(Ɛ��}�l
�O�)��Բ�>o�����ާ�)�u�p�S��>}z����"y�|���꭮�$B�6��mlׇ�.�$v��E' x�^wj\�A1��Rd'�F~	�M���8)���O�s3���0��5�I(MN�#8^e2�y��t�nG���p�}#)Qy���������Mگs�K]s|i�Yg�++�$���IPвP�;=O�mEA�qR�k9g� �)��\B��[�LÑ�D� �փtݻy��'���}���8xknd�W�ff���$^�rD��+kN�7:�����q��;tj�_Շf�'���Lv�n�F�UP>���7
$�ſdIw��	P`�o�,�R{�)��1�14�=�� ����t�*E�EE����Ƽ/��QOc��)1K��zg`i]"�7�PH#�j툞�.�+χ)� UK���Z&j�%ͥ�r���(������Ui��B��~A�[��'�sd��K�zI7�~I�))�V�w�A�2��혏1����ޑ0�"�d,N(|�Jk��3��G6�aG5lZS\��Y[�4%���/���8�R�v^�������(~b��kFrL���>C[�k��,����Q�~�Q�Jj2����\����YQ��Aa�S�zx<4�A�(��k�g��amD��҅tOa���t!�'f^5B������މ����k�ޚ�֑�{p��l4D�.�x� ��LKqߛˈ�ϔnE�Q�ţ�#J[L�>@��NT���F|ڪ�J���){�'��b-��
)�Ԩ�4m�}=L�����P
��	Y�ދ�B�͔[�)�!�9�eU���U�"e���$��+>T�����\j�.G?3ci)��ZDQP��f�V�Ê!�~> (���S��͡�f��r�tU��O� n�Q:
n�s�UЙ��́��#c��d8���Q*(
��C�BG��H��2�k�?Fx���.�k�Ǒw�����5g�Pi�)�մ���\d����@+����	p\:��sε�d�o$�$cn�v2p߂bpGU�|do��Z����|�X�u!W,P^U�._U{��D�B�z�hwᘥHeY	V)w�-a[�����4��M��U�nU��Q�׫����'�J���e�E�+	aU�L	�rO��i$�@��W�ԩb�b�~�V���.(B��ҰY"��U�ժ\����l��/lir��U��&dO���\��eJ��%���?�@H6$Y^
�oW�W�@I(��}Ov���v�R� Ť�$uz�j�#��~�B(�R@!c��T�Ga;��Ps%��Hh:
�y�ݶ�F��1��
|u�����᪒%W�-ۡ ��Z�,���&TFR��[��*��[�Q2�v�*���?ER:�W��0��}��{��)C"�#��}���P?�u�([�ز�����o��� �N0\�d���`��Aβ��f��/RU-��T(2"��44Y
7���d��@>"�
L�|t�x����6�g|�/�$��s](�����#�3��s��4"_rO�OE�$KF���'!��AI2�@;s�����9��Y�R����|��ç�9����qsHD�Z;|���O	��|E�Kd��Z���0
4���S�kE
���Rx-�c��ُ��S(�IRd�쑔���r�Q~� �A�.脳�1(���H�2]�5���?ES���)�y_�.
]x�3~ ��f|�{	)�����|F�}��i��%I��3:����]ܻw��~���q�9��?R܏d+a��%䶾����]Ɠ\�<� ���$�e�(��RD̴A�RD�B�""A@_���6ĎM!��Q�l(08
	�DH�Wǉ8Q)��E��)��$����a!�^!���"2�RD����|��P����ryv*|�
y��q\/-�kE�Y"ŭD&r�t����((
����((
����((
��P���b(@b(HR�w@�R�,����RH!��?Q9����|    IEND�B`�PK   �\XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   �\X ��  u(     jsons/user_defined.json�[o�6ǿ��l�i�N*o��v�$ȭ� �(�jK�,7͊~�ɗđ��m�<Ħ�����\��_=�\������.qi���?�q�<+r����|ח��G�~[85�z�LY^��O��Bk*��(����̖�-�,&W�o�Aǫs�R3��A?��}ʒXp̐#űE�����s�dǱ��2�UK#���3�SN�E��U�	���BJ9�,��5��a_�9�	fyG�Ky���b��'yZ�����8��&�q\L浭�P�%O��C�N��^Z���X��$�U��q����b�Ն��&�B����/��(��E	[�GU� �LL�ꫮO�/���������ؕ��ܓ��7o�X�Ɗ 셛�ʋem�²!��Ry������m�b�;�?,نF?U-(�A�X�AuJ��#�eFm�G/���mYѰ�Q?�-*�#懶%E�b��ж�hX菄��S�ůB/������ۡ)��J��-+Bø��J��",{LvW[[��b�B�EK�b���EK�b���v-���Ԏ����Omk���!T姶5FI U��m�5� ���2��n�@�?!Ҏ���~yю�%�~u���%�~q������ۦ��Z�Y	��w�������I�EV�8�)����w�Sj�MKW��,f����谚7�KC��^��Y^�f�h&
��:��ުU�_<���b:�X\�7�<�'n�V�ϋ�ަ����;����jQ�`���� ��Z�R�.�n��/N�G�ws�rx���ɝ5��5�s{�zsy���=��0�}��f��E��s�g���re�^�����V�qk9R4�VD�$&I��#�5G����q"���&tڒ�"�Kq��0&e������P�
��<68���U�F2Il"I��h�i��v�i�^F|kVSCZ���4r9B#���=�]���ܶ�����W�:����@�n`�Y$�xm����c����RCF%{3�1�Q�k��~��чu�?����O���齣jn�}����k�[�.� ���[	�3��v�Jaw�LL9}���!!���v���S8I��"B,$�@6rYb	'`>���L�.(k�$��,���p&�i�	����d1U̴�,ZM kY,4�I�Q��b�#1�J�?���P�Ku%-��Q�x�?3��� ��PpB^I[;F���B�J��2�s��=T�NZbo~��B�Җ�S������!�v�@�4<�Ȱ(BP���r�!IRc8S��4�dG�]rN�P��E�E)'$�q��dݿmE�yu��yg��2+<9bZ|1u[���N��!�&�r_�^\|���`!;��^U�\�Ul5gކoc��g+��j�w�y��A?�d��:�/?d����ͦg&<��cY,�D^<o8{ۼ��x63v�Ȟ���-�0^5N{��"�.���3c� �2.e%��=�2�v+K�R&:J�BLC�v�N!M��0��Tū���A�=�|��A�=�|��A�=�|��A�=�������PK   �\XL�Q�  yj            ��    cirkitFile.jsonPK   �\XH�8�  �  /           ���  images/273c8146-c058-4dd4-bed5-b60da603675f.pngPK   �\X����7  �  /           ��.  images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK   �\X|�K�?  :  /           ���?  images/54ba0d46-ef45-4902-8525-adba90967d59.pngPK   �\X��@��  ֈ  /           ��U  images/6b718467-4333-41a0-af30-09c4429f5121.pngPK   �\X�&�}[  y`  /           ��}�  images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK   �\X$7h�!  �!  /           ��G2 images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK   �\X�����  �  /           ���T images/edbb92c6-3c2c-4408-8481-9459a63b273a.pngPK   �\XP��/�  ǽ  /           ���k images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK   �\X ��  u(             �� jsons/user_defined.jsonPK    
 
 j  O$   